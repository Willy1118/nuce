module pattern(row_bin, col);

	input [3:0] row_bin;
	output reg [15:0] col;
	
	always @(*) begin
		case(row_bin)
			4'd0:  col = 16'b0000000000000000;
			4'd1:  col = 16'b0000110000000000;
			4'd2:  col = 16'b0001111000000000;
			4'd3:  col = 16'b0000110000000000;
			4'd4:  col = 16'b0000011000000000;
			4'd5:  col = 16'b0000011110000000;
			4'd6:  col = 16'b0000011101000000;
			4'd7:  col = 16'b0000101101000000;
			4'd8:  col = 16'b0001001100000000;
			4'd9:  col = 16'b0000001110000000;
			4'd10: col = 16'b0000001010000000;
			4'd11: col = 16'b0000010001100000;
			4'd12: col = 16'b0000010000011000;
			4'd13: col = 16'b0000010000001000;
			4'd14: col = 16'b0001100000010000;
			4'd15: col = 16'b0000000000000000;
			default: col = 16'b0000000000000000;
		endcase
	end

endmodule 